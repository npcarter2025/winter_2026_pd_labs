
.SUBCKT INVx4_ASAP7_6t_R A VDD VSS Y
MM0 Y A VSS VSS nmos_rvt w=216.00n l=20n nfin=8
MM1 Y A VDD VDD pmos_rvt w=216.00n l=20n nfin=8
.ENDS